/*
DVI Test Top Module
retrocpu DVI Character Display GPU - Phase 3 Hardware Validation

Top-level module for validating DVI output with test patterns.
Integrates:
- PLL (25 MHz → 125 MHz TMDS clock + 25 MHz pixel clock)
- VGA timing generator (640x480@60Hz)
- Test pattern generator
- DVI transmitter with TMDS encoding
- ECP5 LVDS output primitives

Target: Colorlight i5 v7.0
Created: 2025-12-28
*/

module dvi_test_top(
    input  wire       clk_25mhz,      // 25 MHz oscillator input

    output wire [3:0] gpdi_dp,        // TMDS data positive (3=clk, 2=red, 1=green, 0=blue)
    // Note: gpdi_dn is not declared - LVCMOS33D mode automatically generates differential negative signals

    output wire       led             // Status LED (blinks at frame rate)
);

// Test pattern selection (hardcoded for now)
// 00 = Color bars, 01 = Checkerboard, 10 = Grid, 11 = Solid gray
wire [1:0] pattern_sel = 2'b00;  // Color bars pattern

//=============================================================================
// Clock Generation (PLL)
//=============================================================================

wire [3:0] clocks;
wire       pll_locked;

ecp5_pll #(
    .in_hz(25_000_000),      // 25 MHz input
    .out0_hz(125_000_000),   // TMDS clock (5x pixel clock for DDR)
    .out1_hz(25_000_000)     // Pixel clock
) pll_inst (
    .clk_i(clk_25mhz),
    .clk_o(clocks),
    .locked(pll_locked),
    // Tie off unused ports
    .reset(1'b0),
    .standby(1'b0),
    .phasesel(2'b00),
    .phasedir(1'b0),
    .phasestep(1'b0),
    .phaseloadreg(1'b0)
);

wire tmds_clk = clocks[0];  // 125 MHz
wire pclk     = clocks[1];  // 25 MHz

// Generate reset from PLL lock
reg [3:0] reset_count = 0;
reg rst_n = 0;

always @(posedge pclk) begin
    if (pll_locked) begin
        if (reset_count != 4'hF) begin
            reset_count <= reset_count + 1;
        end else begin
            rst_n <= 1;
        end
    end else begin
        reset_count <= 0;
        rst_n <= 0;
    end
end

//=============================================================================
// VGA Timing Generator (using reference implementation)
//=============================================================================

wire [10:0] h_count;
wire [10:0] v_count;
wire       hsync;
wire       vsync;
wire       blank;

my_vga_clk_generator vga_timing_inst (
    .pclk(pclk),
    .reset_n(rst_n),
    .out_hcnt(h_count),
    .out_vcnt(v_count),
    .out_hsync(hsync),
    .out_vsync(vsync),
    .out_blank(blank)
);

// Derive video_active and frame_start
wire video_active = ~blank;
wire frame_start = (h_count == 0) && (v_count == 0);

//=============================================================================
// Test Pattern Generator
//=============================================================================

wire [7:0] red;
wire [7:0] green;
wire [7:0] blue;

test_pattern_generator test_pattern_inst (
    .clk(pclk),
    .rst_n(rst_n),
    .h_count(h_count),
    .v_count(v_count),
    .video_active(video_active),
    .pattern_sel(pattern_sel),
    .red(red),
    .green(green),
    .blue(blue)
);

//=============================================================================
// DVI Transmitter (TMDS Encoding + Serialization)
//=============================================================================

wire [1:0] tmds_red;
wire [1:0] tmds_green;
wire [1:0] tmds_blue;
wire [1:0] tmds_clock;

dvi_transmitter dvi_transmitter_inst (
    .pclk(pclk),
    .tmds_clk(tmds_clk),
    .in_red(red),
    .in_green(green),
    .in_blue(blue),
    .in_blank(~video_active),
    .in_vsync(vsync),
    .in_hsync(hsync),
    .out_tmds_red(tmds_red),
    .out_tmds_green(tmds_green),
    .out_tmds_blue(tmds_blue),
    .out_tmds_clk(tmds_clock)
);

//=============================================================================
// ECP5 LVDS Output Primitives (DDR)
//=============================================================================

// TMDS Clock output
ODDRX1F ddr_clk (
    .D0(tmds_clock[0]),
    .D1(tmds_clock[1]),
    .Q(gpdi_dp[3]),
    .SCLK(tmds_clk),
    .RST(1'b0)
);

// TMDS Red output
ODDRX1F ddr_red (
    .D0(tmds_red[0]),
    .D1(tmds_red[1]),
    .Q(gpdi_dp[2]),
    .SCLK(tmds_clk),
    .RST(1'b0)
);

// TMDS Green output
ODDRX1F ddr_green (
    .D0(tmds_green[0]),
    .D1(tmds_green[1]),
    .Q(gpdi_dp[1]),
    .SCLK(tmds_clk),
    .RST(1'b0)
);

// TMDS Blue output
ODDRX1F ddr_blue (
    .D0(tmds_blue[0]),
    .D1(tmds_blue[1]),
    .Q(gpdi_dp[0]),
    .SCLK(tmds_clk),
    .RST(1'b0)
);

// Note: gpdi_dn outputs are automatically generated by LVCMOS33D IO type
// (differential mode in the LPF file - no explicit assignment needed)

//=============================================================================
// Status LED (frame rate indicator)
//=============================================================================

// Blink LED at ~1Hz (count 60 frames)
reg [5:0] frame_count = 0;
reg led_state = 0;

always @(posedge pclk) begin
    if (frame_start) begin
        if (frame_count == 59) begin
            frame_count <= 0;
            led_state <= ~led_state;
        end else begin
            frame_count <= frame_count + 1;
        end
    end
end

assign led = led_state;

endmodule
